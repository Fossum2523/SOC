// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module exmem #(
    parameter BITS = 32,
    parameter DELAYS=10
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wire wbs_clk_i,
    input wire wbs_rst_i,
    input wire [31:0] wbs_adr_i,
    input wire [31:0] wbs_dat_i,
    input wire [3:0] wbs_sel_i,
    input wire wbs_we_i,
    input wire wbs_cyc_i,
    input wire wbs_stb_i,
    input wire wbs_err_i,
    output reg wbs_ack_o,
    output wire [31:0] wbs_dat_o

    // Logic Analyzer Signals
   /* input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq*/
);
    wire clk;
    wire rst;

    /*wire [`MPRJ_IO_PADS-1:0] io_in;
    wire [`MPRJ_IO_PADS-1:0] io_out;
    wire [`MPRJ_IO_PADS-1:0] io_oeb;*/
    wire [31:0]addr;
    wire decode;
    wire [31:0]data_out;
    wire EN0;
    wire [3:0]wstrb;
    
    assign clk = wbs_clk_i;
    assign rst = wbs_rst_i;
    //assign addr = wbs_adr_i - 32'h38000000;
    assign decode = wbs_adr_i[31:20] == 12'h380 ? 1'b1:1'b0;
    assign wbs_dat_o = (wbs_ack_o) ?data_out:32'd0;
    assign EN0 = wbs_stb_i && wbs_cyc_i && decode;
    //assign wbs_dat_o = 32'd0;
    assign wstrb = wbs_sel_i &{4{wbs_we_i}};
    
    bram user_bram (
        .CLK(clk),
        .WE0(wstrb),
        .EN0(EN0),
        .Di0(wbs_dat_i),
        .Do0(data_out),
        .A0(wbs_adr_i)
        //.A0(addr)
    );
    
    reg [3:0]counter;
    
    always @(posedge clk)begin
    	if(rst)begin	
    	   counter <= 4'd0;
    	   wbs_ack_o <= 1'd0;
    	end
    	else begin
    	   if(wbs_stb_i && wbs_cyc_i)begin
    	   	
    	   	if(counter==DELAYS)begin
    	   	    wbs_ack_o <= 1'd1;
    	   	    
    	   	    counter <= 4'd0;
    	   	end
    	   	else begin
    	   	    counter <= counter + 4'd1;
    	   	    wbs_ack_o <= 1'd0;
    	   	end
    	   end
    	   else begin
    	   	counter <= 4'd0;
    	   	
    	   end
    	end
    end
	
	
	
endmodule



`default_nettype wire